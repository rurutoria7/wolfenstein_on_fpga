module Raycaster;
endmodule;